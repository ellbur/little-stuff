
Vs 1 0 pulse(0 5 0 0 0 0.5ms 1ms)
R1 1 0 10k

.tran 0.01ms 2ms

