
.subckt src p n
V p n PWL(
+ 0.0 0.0
+ 0.0 1.0
+ 0.0204081632653 0.991790013823
+ 0.0408163265306 0.967294863039
+ 0.0612244897959 0.926916757346
+ 0.0816326530612 0.871318704123
+ 0.102040816327 0.801413621868
+ 0.122448979592 0.718349350098
+ 0.142857142857 0.623489801859
+ 0.163265306122 0.518392568311
+ 0.183673469388 0.404783343122
+ 0.204081632653 0.284527586631
+ 0.224489795918 0.159599895033
+ 0.244897959184 0.0320515775717
+ 0.265306122449 -0.0960230259077
+ 0.285714285714 -0.222520933956
+ 0.30612244898 -0.345365054421
+ 0.326530612245 -0.462538290241
+ 0.34693877551 -0.572116660122
+ 0.367346938776 -0.672300890261
+ 0.387755102041 -0.761445958369
+ 0.408163265306 -0.838088104892
+ 0.428571428571 -0.900968867902
+ 0.448979591837 -0.949055747011
+ 0.469387755102 -0.981559156991
+ 0.489795918367 -0.99794539275
+ 0.510204081633 -0.99794539275
+ 0.530612244898 -0.981559156991
+ 0.551020408163 -0.949055747011
+ 0.571428571429 -0.900968867902
+ 0.591836734694 -0.838088104892
+ 0.612244897959 -0.761445958369
+ 0.632653061224 -0.672300890261
+ 0.65306122449 -0.572116660122
+ 0.673469387755 -0.462538290241
+ 0.69387755102 -0.345365054421
+ 0.714285714286 -0.222520933956
+ 0.734693877551 -0.0960230259077
+ 0.755102040816 0.0320515775717
+ 0.775510204082 0.159599895033
+ 0.795918367347 0.284527586631
+ 0.816326530612 0.404783343122
+ 0.836734693878 0.518392568311
+ 0.857142857143 0.623489801859
+ 0.877551020408 0.718349350098
+ 0.897959183673 0.801413621868
+ 0.918367346939 0.871318704123
+ 0.938775510204 0.926916757346
+ 0.959183673469 0.967294863039
+ 0.979591836735 0.991790013823
+ 1.0 1.0
+ 1.0 1.0
+ 1.02040816327 0.967294863039
+ 1.04081632653 0.871318704123
+ 1.0612244898 0.718349350098
+ 1.08163265306 0.518392568311
+ 1.10204081633 0.284527586631
+ 1.12244897959 0.0320515775717
+ 1.14285714286 -0.222520933956
+ 1.16326530612 -0.462538290241
+ 1.18367346939 -0.672300890261
+ 1.20408163265 -0.838088104892
+ 1.22448979592 -0.949055747011
+ 1.24489795918 -0.99794539275
+ 1.26530612245 -0.981559156991
+ 1.28571428571 -0.900968867902
+ 1.30612244898 -0.761445958369
+ 1.32653061224 -0.572116660122
+ 1.34693877551 -0.345365054421
+ 1.36734693878 -0.0960230259077
+ 1.38775510204 0.159599895033
+ 1.40816326531 0.404783343122
+ 1.42857142857 0.623489801859
+ 1.44897959184 0.801413621868
+ 1.4693877551 0.926916757346
+ 1.48979591837 0.991790013823
+ 1.51020408163 0.991790013823
+ 1.5306122449 0.926916757346
+ 1.55102040816 0.801413621868
+ 1.57142857143 0.623489801859
+ 1.59183673469 0.404783343122
+ 1.61224489796 0.159599895033
+ 1.63265306122 -0.0960230259077
+ 1.65306122449 -0.345365054421
+ 1.67346938776 -0.572116660122
+ 1.69387755102 -0.761445958369
+ 1.71428571429 -0.900968867902
+ 1.73469387755 -0.981559156991
+ 1.75510204082 -0.99794539275
+ 1.77551020408 -0.949055747011
+ 1.79591836735 -0.838088104892
+ 1.81632653061 -0.672300890261
+ 1.83673469388 -0.462538290241
+ 1.85714285714 -0.222520933956
+ 1.87755102041 0.0320515775717
+ 1.89795918367 0.284527586631
+ 1.91836734694 0.518392568311
+ 1.9387755102 0.718349350098
+ 1.95918367347 0.871318704123
+ 1.97959183673 0.967294863039
+ 2.0 1.0
+ 2.0 1.0
+ 2.02040816327 0.926916757346
+ 2.04081632653 0.718349350098
+ 2.0612244898 0.404783343122
+ 2.08163265306 0.0320515775717
+ 2.10204081633 -0.345365054421
+ 2.12244897959 -0.672300890261
+ 2.14285714286 -0.900968867902
+ 2.16326530612 -0.99794539275
+ 2.18367346939 -0.949055747011
+ 2.20408163265 -0.761445958369
+ 2.22448979592 -0.462538290241
+ 2.24489795918 -0.0960230259077
+ 2.26530612245 0.284527586631
+ 2.28571428571 0.623489801859
+ 2.30612244898 0.871318704123
+ 2.32653061224 0.991790013823
+ 2.34693877551 0.967294863039
+ 2.36734693878 0.801413621868
+ 2.38775510204 0.518392568311
+ 2.40816326531 0.159599895033
+ 2.42857142857 -0.222520933956
+ 2.44897959184 -0.572116660122
+ 2.4693877551 -0.838088104892
+ 2.48979591837 -0.981559156991
+ 2.51020408163 -0.981559156991
+ 2.5306122449 -0.838088104892
+ 2.55102040816 -0.572116660122
+ 2.57142857143 -0.222520933956
+ 2.59183673469 0.159599895033
+ 2.61224489796 0.518392568311
+ 2.63265306122 0.801413621868
+ 2.65306122449 0.967294863039
+ 2.67346938776 0.991790013823
+ 2.69387755102 0.871318704123
+ 2.71428571429 0.623489801859
+ 2.73469387755 0.284527586631
+ 2.75510204082 -0.0960230259077
+ 2.77551020408 -0.462538290241
+ 2.79591836735 -0.761445958369
+ 2.81632653061 -0.949055747011
+ 2.83673469388 -0.99794539275
+ 2.85714285714 -0.900968867902
+ 2.87755102041 -0.672300890261
+ 2.89795918367 -0.345365054421
+ 2.91836734694 0.0320515775717
+ 2.9387755102 0.404783343122
+ 2.95918367347 0.718349350098
+ 2.97959183673 0.926916757346
+ 3.0 1.0
+ 3.0 1.0
+ 3.02040816327 0.871318704123
+ 3.04081632653 0.518392568311
+ 3.0612244898 0.0320515775717
+ 3.08163265306 -0.462538290241
+ 3.10204081633 -0.838088104892
+ 3.12244897959 -0.99794539275
+ 3.14285714286 -0.900968867902
+ 3.16326530612 -0.572116660122
+ 3.18367346939 -0.0960230259077
+ 3.20408163265 0.404783343122
+ 3.22448979592 0.801413621868
+ 3.24489795918 0.991790013823
+ 3.26530612245 0.926916757346
+ 3.28571428571 0.623489801859
+ 3.30612244898 0.159599895033
+ 3.32653061224 -0.345365054421
+ 3.34693877551 -0.761445958369
+ 3.36734693878 -0.981559156991
+ 3.38775510204 -0.949055747011
+ 3.40816326531 -0.672300890261
+ 3.42857142857 -0.222520933956
+ 3.44897959184 0.284527586631
+ 3.4693877551 0.718349350098
+ 3.48979591837 0.967294863039
+ 3.51020408163 0.967294863039
+ 3.5306122449 0.718349350098
+ 3.55102040816 0.284527586631
+ 3.57142857143 -0.222520933956
+ 3.59183673469 -0.672300890261
+ 3.61224489796 -0.949055747011
+ 3.63265306122 -0.981559156991
+ 3.65306122449 -0.761445958369
+ 3.67346938776 -0.345365054421
+ 3.69387755102 0.159599895033
+ 3.71428571429 0.623489801859
+ 3.73469387755 0.926916757346
+ 3.75510204082 0.991790013823
+ 3.77551020408 0.801413621868
+ 3.79591836735 0.404783343122
+ 3.81632653061 -0.0960230259077
+ 3.83673469388 -0.572116660122
+ 3.85714285714 -0.900968867902
+ 3.87755102041 -0.99794539275
+ 3.89795918367 -0.838088104892
+ 3.91836734694 -0.462538290241
+ 3.9387755102 0.0320515775716
+ 3.95918367347 0.518392568311
+ 3.97959183673 0.871318704123
+ 4.0 1.0
+ )
.ends

