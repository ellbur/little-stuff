
.include source.sp

X1 1 0 src
R1 1 0 1k

.tran 0.01, 4

